module spi_MBslave(
    input clk,
    input rst,
    input ss,
    input mosi,
    output miso,
    input sck,
    output done,
    input [7:0] din,
    output [7:0] dout
    );

//parameter buffersize 



//spi_slave spi_slave (clk, rst, ss, mosi,miso,sck, done, din, dout);

endmodule
